module ghost()